
/******************************************************************************
 Copyright (c) 2004-2018, AMIQ Consulting srl. All rights reserved.

 Licensed under the Apache License, Version 2.0 (the "License");
 you may not use this file except in compliance with the License.
 You may obtain a copy of the License at
 http://www.apache.org/licenses/LICENSE-2.0

 Unless required by applicable law or agreed to in writing, software
 distributed under the License is distributed on an "AS IS" BASIS,
 WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 See the License for the specific language governing permissions and
 limitations under the License.
 *******************************************************************************/

`ifndef __EX_ENV
`define __EX_ENV

class ex_env extends uvm_env;
	`uvm_component_utils(ex_env)
	// Components of the environment
	//TODO: instantiate here
	ex_in_agent in_agent;
	ex_out_agent out_agent;
	ex_scoreboard sb;

	function new(string name, uvm_component parent);
		super.new(name, parent);
	endfunction : new

	virtual function void build_phase(uvm_phase phase);
		super.build_phase(phase);
		//TODO: create agents and others here
		in_agent  = ex_in_agent::type_id::create(.name("in_agent"), .parent(this));
		in_agent.is_active = UVM_ACTIVE;
		out_agent  = ex_out_agent::type_id::create(.name("out_agent"), .parent(this));
		sb = ex_scoreboard::type_id::create("scoreboard", this);
	endfunction : build_phase

	function void connect_phase (uvm_phase phase);
		//TODO: connect stuff here
		super.connect_phase(phase);      
		in_agent.monitor.collected_item_port.connect(sb.in_port);      
		out_agent.monitor.collected_item_port.connect(sb.out_port);
	endfunction : connect_phase

endclass : ex_env

`endif



